module cpu (clk, reset, instruction, data_out);
input clk;
input reset;
input [7:0] instruction;
output reg [7:0] data_out;

//register declaration

//ALU?

//control unit

//pc (program counter)

//data memory

//instruction memory

always @(*) begin
    //top
end

endmodule